interface alu_interface(input logic clk); 
  
  logic in;
  logic out;
  logic sign;
  logic carr;
  logic zero;
  
endinterface:alu_interface